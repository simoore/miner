///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module MinerCore(
    input logic clk
);
    
    Hasher hasher0 (
    );
    
    
endmodule



