package Sha256Types;



endpackage