import Sha256Types::*;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module MinerCore(

    );
    
    
    
endmodule



