module MinerTop (

);

endmodule
