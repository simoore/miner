package Sha256Types;

typedef logic [31:0] uint32_t;

typedef struct {
    uint32_t a;
    uint32_t b;
    uint32_t c;
    uint32_t d;
    uint32_t e;
    uint32_t f;
    uint32_t g;
    uint32_t h;
} WorkingVars;

endpackage